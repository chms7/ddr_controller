// module mc_dfi_if #(
//   parameter FREQ_RAT_PHY2MC = 4;
// ) (

// );
  
// endmodule
